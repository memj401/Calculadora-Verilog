module pilha( 
    input  tecla[3:0],
	 output [4:0] A,
	 output [4:0] B,
    );